/home/ashish/FileSystemTest/Sem4/COL216/2017CS10389_2017CS50521/Testbench.vhd